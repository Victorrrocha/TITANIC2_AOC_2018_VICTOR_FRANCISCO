LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RAM16 IS
PORT(
	CLOCK	: 	IN 	STD_LOGIC;
	ROW	: 	IN 	STD_LOGIC; 								--READ OR WRITE
	ADDRESS:	IN 	STD_LOGIC_VECTOR (3 DOWNTO 0); 	--ENDEREÇO PARA ROW
	DATAIN:	IN 	STD_LOGIC_VECTOR (15 DOWNTO 0); 	--DADO A SER ESCRITO
	DATAOUT:	OUT	STD_LOGIC_VECTOR (15 DOWNTO 0) 	--DADO A SER LIDO
);
END ENTITY RAM16;

ARCHITECTURE RAM_BH OF RAM16 IS

	TYPE RAM_ARRAY IS ARRAY (15 DOWNTO 0)  OF STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL RAM : RAM_ARRAY; -- instanciando uma estrutura ram_bh
	SIGNAL READ_ADDRESS : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN 
	PROCESS(CLOCK) IS
	
	BEGIN
		IF RISING_EDGE(CLOCK) THEN
			IF ROW = '0' THEN --ARMAZENANDO
				RAM(TO_INTEGER(UNSIGNED(ADDRESS))) <= DATAIN;
			END IF;
			READ_ADDRESS <= ADDRESS;
		END IF;
	END PROCESS;
	
	DATAOUT <= RAM(TO_INTEGER(UNSIGNED(READ_ADDRESS))) WHEN ROW = '1';

END ARCHITECTURE RAM_BH;